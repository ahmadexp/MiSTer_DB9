//=========================================================
//  Arcade: SEGA SYSTEM 1  for MiSTer
//
//                          Copyright (c) 2019 MiSTer-X
//=========================================================

module emu
(
	//Master input clock
	input         CLK_50M,

	//Async reset from top-level module.
	//Can be used as initial reset.
	input         RESET,

	//Must be passed to hps_io module
	inout  [45:0] HPS_BUS,

	//Base video clock. Usually equals to CLK_SYS.
	output        VGA_CLK,

	//Multiple resolutions are supported using different VGA_CE rates.
	//Must be based on CLK_VIDEO
	output        VGA_CE,

	output  [7:0] VGA_R,
	output  [7:0] VGA_G,
	output  [7:0] VGA_B,
	output        VGA_HS,
	output        VGA_VS,
	output        VGA_DE,    // = ~(VBlank | HBlank)
	output		  VGA_F1,
	
	//Base video clock. Usually equals to CLK_SYS.
	output        HDMI_CLK,

	//Multiple resolutions are supported using different HDMI_CE rates.
	//Must be based on CLK_VIDEO
	output        HDMI_CE,

	output  [7:0] HDMI_R,
	output  [7:0] HDMI_G,
	output  [7:0] HDMI_B,
	output        HDMI_HS,
	output        HDMI_VS,
	output        HDMI_DE,   // = ~(VBlank | HBlank)
	output  [1:0] HDMI_SL,   // scanlines fx

	//Video aspect ratio for HDMI. Most retro systems have ratio 4:3.
	output  [7:0] HDMI_ARX,
	output  [7:0] HDMI_ARY,
	
	//DB9 Joystick
	input [5:0] joy_o_db9,    // CB UDLR
	output      db9_Select,
	output      splitter_select,
	
	output        LED_USER,  // 1 - ON, 0 - OFF.

	// b[1]: 0 - LED status is system status OR'd with b[0]
	//       1 - LED status is controled solely by b[0]
	// hint: supply 2'b00 to let the system control the LED.
	output  [1:0] LED_POWER,
	output  [1:0] LED_DISK,

	output [15:0] AUDIO_L,
	output [15:0] AUDIO_R,
	output        AUDIO_S,   // 1 - signed audio samples, 0 - unsigned

	// Open-drain User port.
	// 0 - D+/RX
	// 1 - D-/TX
	// 2..6 - USR2..USR6
	// Set USER_OUT to 1 to read from USER_IN.
	input   [6:0] USER_IN,
	output  [6:0] USER_OUT
);

assign VGA_F1    = 0;
assign USER_OUT  = '1;
assign LED_USER  = ioctl_download;
assign LED_DISK  = 0;
assign LED_POWER = 0;

wire   screen_H = status[6]|~SYSMODE[1]|direct_video;
assign HDMI_ARX = status[1] ? 8'd16 : screen_H ? 8'd4 : 8'd3;
assign HDMI_ARY = status[1] ? 8'd9  : screen_H ? 8'd3 : 8'd4;

`include "build_id.v" 

localparam CONF_STR = {
	"A.SEGASYS1;;",
	"-;",
	"H0O1,Aspect Ratio,Original,Wide;",
	"O35,Scandoubler Fx,None,HQ2x,CRT 25%,CRT 50%,CRT 75%;",
	"H0O6,Auto Rotation,On,Off;",
	"-;",
	"DIP;",
	"-;",
	"OOS,Analog Video H-Pos,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30,31;",
	"OTV,Analog Video V-Pos,0,1,2,3,4,5,6,7;",
	"-;",
	"R0,Reset;",
	"J1,Trig1,Trig2,Trig3,Start 1P,Start 2P,Coin;",
	"jn,A,B,R,Start,Select,L;",
	"V,v",`BUILD_DATE
};

wire bCabinet = 1'b0;

wire [4:0] HOFFS = status[28:24];
wire [2:0] VOFFS = status[31:29];

//////  I/O TWO JOYSTICK SPLITTER OPTION ADDED FROM JOYAV //////////

//assign db9_Select = 1'b1;
assign splitter_select = 1'bz; 
wire [5:0] JOYAV_T1;      // CB UDLR  negative Logic

assign JOYAV_T1 = joy_o_db9; 

// Now we apply the megadrive desmultiplexor conversor
wire [11:0] joy1_o;   // MXYZ SACB RLDU  in negative logic

// Then, we call the states machine to read the six Megadrive controller buttons
// Format joy1_o [11:0] =  MXYZ SACB RLDU negative logic
sega_joystick joy_megadrive (
	.joy1_up_i		(JOYAV_T1[3]), // JOYAV_T1 // CB UDLR (negative logic)
	.joy1_down_i	(JOYAV_T1[2]),
	.joy1_left_i	(JOYAV_T1[1]),
	.joy1_right_i	(JOYAV_T1[0]),
	.joy1_p6_i		(JOYAV_T1[4]),
	.joy1_p9_i		(JOYAV_T1[5]),
	.vga_hsync_n_s (hblank),
	.joyX_p7_o		(db9_Select), // select signal
	.joy1_o			(joy1_o)    // MXYZ SACB RLDU in negative logic
); 
							// Coin,    Start 2P,    Start 1P,     T3, 			T2, 			T1,  		   RLDU
wire [9:0] JOYAV_1;  //  M           Z           S           A      		 B     		C			   UDLR   in positive logic

assign JOYAV_1 = ~{ joy1_o[11],   joy1_o[8],   joy1_o[7], joy1_o[6],	 joy1_o[5],  joy1_o[4],   joy1_o[0],joy1_o[1],joy1_o[2],joy1_o[3]};  



////////////////////   CLOCKS   ///////////////////

wire clk_48M;
wire clk_hdmi = clk_48M;
wire clk_sys  = clk_48M;

pll pll
(
	.rst(0),
	.refclk(CLK_50M),
	.outclk_0(clk_48M)
);

///////////////////////////////////////////////////

wire [31:0] status;
wire  [1:0] buttons;
wire        forced_scandoubler;
wire			direct_video;

wire        ioctl_download;
wire        ioctl_wr;
wire  [7:0]	ioctl_index;
wire [24:0] ioctl_addr;
wire  [7:0] ioctl_dout;

wire [10:0] ps2_key;
wire [15:0] joystk1, joystk2;
wire [15:0] joystick_analog_0;
wire [15:0] joystick_analog_1;

wire [21:0]	gamma_bus;

hps_io #(.STRLEN($size(CONF_STR)>>3)) hps_io
(
	.clk_sys(clk_sys),
	.HPS_BUS(HPS_BUS),

	.conf_str(CONF_STR),

	.buttons(buttons),

	.status(status),
	.status_menumask({15'h0,direct_video}),
	
	.forced_scandoubler(forced_scandoubler),
	.gamma_bus(gamma_bus),
	.direct_video(direct_video),

	.ioctl_download(ioctl_download),
	.ioctl_wr(ioctl_wr),
	.ioctl_addr(ioctl_addr),
	.ioctl_dout(ioctl_dout),
	.ioctl_index(ioctl_index),

	.joystick_0(joystk1),
	.joystick_1(joystk2),
	.joystick_analog_0(joystick_analog_0),
	.joystick_analog_1(joystick_analog_1),	

	.ps2_key(ps2_key)
);

reg [7:0] SYSMODE;	// [0]=SYS1/SYS2,[1]=H/V,[2]=H256/H240
reg [7:0] DSW[8];
always @(posedge clk_sys) begin
	if (ioctl_wr) begin
		if ((ioctl_index==1  ) && (ioctl_addr==0))   SYSMODE <= ioctl_dout;
		if ((ioctl_index==254) && !ioctl_addr[24:3]) DSW[ioctl_addr[2:0]] <= ioctl_dout;
	end
end

wire       pressed = ps2_key[9];
wire [8:0] code    = ps2_key[8:0];
always @(posedge clk_sys) begin
	reg old_state;
	old_state <= ps2_key[10];
	
	if(old_state != ps2_key[10]) begin
		casex(code)
			'hX75: btn_up          <= pressed; // up
			'hX72: btn_down        <= pressed; // down
			'hX6B: btn_left        <= pressed; // left
			'hX74: btn_right       <= pressed; // right
			'h029: btn_trig1       <= pressed; // space
			'h014: btn_trig2       <= pressed; // ctrl
			'h011: btn_trig3		  <= pressed; // alt
			'h005: btn_one_player  <= pressed; // F1
			'h006: btn_two_players <= pressed; // F2

			// JPAC/IPAC/MAME Style Codes
			'h016: btn_start_1     <= pressed; // 1
			'h01E: btn_start_2     <= pressed; // 2
			'h02E: btn_coin_1      <= pressed; // 5
			'h036: btn_coin_2      <= pressed; // 6
			'h02D: btn_up_2        <= pressed; // R
			'h02B: btn_down_2      <= pressed; // F
			'h023: btn_left_2      <= pressed; // D
			'h034: btn_right_2     <= pressed; // G
			'h01C: btn_trig1_2     <= pressed; // A
			'h01B: btn_trig2_2     <= pressed; // S
			'h015: btn_trig3_2     <= pressed; // Q
		endcase
	end
end

reg btn_up    = 0;
reg btn_down  = 0;
reg btn_right = 0;
reg btn_left  = 0;
reg btn_trig1 = 0;
reg btn_trig2 = 0;
reg btn_trig3 = 0;
reg btn_one_player  = 0;
reg btn_two_players = 0;

reg btn_start_1 = 0;
reg btn_start_2 = 0;
reg btn_coin_1  = 0;
reg btn_coin_2  = 0;
reg btn_up_2    = 0;
reg btn_down_2  = 0;
reg btn_left_2  = 0;
reg btn_right_2 = 0;
reg btn_trig1_2 = 0;
reg btn_trig2_2 = 0;
reg btn_trig3_2 = 0;



wire m_up2     = btn_up_2    | joystk2[3] | JOYAV_1[3];
wire m_down2   = btn_down_2  | joystk2[2] | JOYAV_1[2];
wire m_left2   = btn_left_2  | joystk2[1] | JOYAV_1[1];
wire m_right2  = btn_right_2 | joystk2[0] | JOYAV_1[0];
wire m_trig21  = btn_trig1_2 | joystk2[4] | JOYAV_1[4];
wire m_trig22  = btn_trig2_2 | joystk2[5] | JOYAV_1[5];
wire m_trig23  = btn_trig3_2 | joystk2[6] | JOYAV_1[6];

wire m_start1  = btn_one_player  | joystk1[7] | joystk2[7] | btn_start_1 | JOYAV_1[7];
wire m_start2  = btn_two_players | joystk1[8] | joystk2[8] | btn_start_2 | JOYAV_1[8];

wire m_up1     = btn_up      | joystk1[3] | (bCabinet ? 1'b0 : m_up2) | JOYAV_1[3];
wire m_down1   = btn_down    | joystk1[2] | (bCabinet ? 1'b0 : m_down2) | JOYAV_1[2];
wire m_left1   = btn_left    | joystk1[1] | (bCabinet ? 1'b0 : m_left2) | JOYAV_1[1];
wire m_right1  = btn_right   | joystk1[0] | (bCabinet ? 1'b0 : m_right2) | JOYAV_1[0];
wire m_trig11  = btn_trig1   | joystk1[4] | (bCabinet ? 1'b0 : m_trig21) | JOYAV_1[4];
wire m_trig12  = btn_trig2   | joystk1[5] | (bCabinet ? 1'b0 : m_trig22) | JOYAV_1[5];
wire m_trig13  = btn_trig3   | joystk1[6] | (bCabinet ? 1'b0 : m_trig23) | JOYAV_1[6];

wire m_coin1   = btn_one_player | btn_coin_1 | joystk1[9] | JOYAV_1[9];
wire m_coin2   = btn_two_players| btn_coin_2 | joystk2[9] | JOYAV_1[9];
wire m_coin    = (m_coin1|m_coin2);


///////////////////////////////////////////////////

wire hblank, vblank;
wire ce_vid;
wire hs, vs;
wire [2:0] r,g;
wire [1:0] b;

reg ce_pix;
always @(posedge clk_hdmi) begin
	reg old_clk;
	old_clk <= ce_vid;
	ce_pix  <= old_clk & ~ce_vid;
end

arcade_rotate_fx #(256,224,8,1) videoV
(
	.*,

	.clk_video(clk_hdmi),

	.RGB_in({r,g,b}),
	.HBlank(hblank),
	.VBlank(vblank),
	.HSync(~hs),
	.VSync(~vs),

	.fx(status[5:3]),
	.no_rotate(screen_H),
);

wire			PCLK;
wire  [8:0] HPOS,VPOS;
wire  [7:0] POUT;
HVGEN hvgen
(
	.HPOS(HPOS),.VPOS(VPOS),.PCLK(PCLK),.iRGB(POUT),
	.oRGB({b,g,r}),.HBLK(hblank),.VBLK(vblank),.HSYN(hs),.VSYN(vs),
	.H240(SYSMODE[2]),.HOFFS(HOFFS),.VOFFS(VOFFS)
);
assign ce_vid = PCLK;


wire [15:0] AOUT;
assign AUDIO_L = AOUT;
assign AUDIO_R = AUDIO_L;
assign AUDIO_S = 0; // unsigned PCM


///////////////////////////////////////////////////

wire iRST = RESET | status[0] | buttons[1];

wire [7:0] INP0 = ~{m_left1,m_right1,m_up1,m_down1,1'd0,m_trig12,m_trig11,m_trig13};
wire [7:0] INP1 = ~{m_left2,m_right2,m_up2,m_down2,1'd0,m_trig22,m_trig21,m_trig23};
wire [7:0] INP2 = ~{2'd0,m_start2,m_start1,3'd0, m_coin}; 


SEGASYSTEM1 GameCore ( 
	.clk48M(clk_48M),.reset(iRST),

	.INP0(INP0),.INP1(INP1),.INP2(INP2),
	.DSW0(DSW[0]),.DSW1(DSW[1]),

	.PH(HPOS),.PV(VPOS),.PCLK(PCLK),.POUT(POUT),
	.SOUT(AOUT),

	.ROMCL(clk_sys),.ROMAD(ioctl_addr),.ROMDT(ioctl_dout),.ROMEN(ioctl_wr & (ioctl_index==0))
);

endmodule

